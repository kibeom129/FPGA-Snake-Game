library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use std.textio.all;

entity random_gen is
  port(
	clk : in std_logic;
  );
end random_gen;

architecture synth of random_gen is

end synth;